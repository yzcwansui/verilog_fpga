
module and_gate
(
a, b, f
);

input a;
input b;
output f;
assign f=a&b;
endmodule
